module test(in,out);
input[31:0] in;
output[9:0] out;

assign out = in[0:9];

endmodule
